module multiplexer (

);


endmodule